library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
library GhdlLink;
use GhdlLink.Utility_Package.all;
use GhdlLink.Vhpi_Foreign.all;
entity ahir_system_Test_Bench is -- 
  -- 
end entity;
architecture VhpiLink of ahir_system_Test_Bench is -- 
  component ahir_system is -- 
    port (-- 
      pmul19_P1 : in  std_logic_vector(15 downto 0);
      pmul19_P2 : in  std_logic_vector(15 downto 0);
      pmul19_result : out  std_logic_vector(15 downto 0);
      pmul19_tag_in: in std_logic_vector(1 downto 0);
      pmul19_tag_out: out std_logic_vector(1 downto 0);
      pmul19_start_req : in std_logic;
      pmul19_start_ack : out std_logic;
      pmul19_fin_req   : in std_logic;
      pmul19_fin_ack   : out std_logic;
      clk : in std_logic;
      reset : in std_logic); -- 
    -- 
  end component;
  signal clk: std_logic := '0';
  signal reset: std_logic := '1';
  signal pmul19_P1 :  std_logic_vector(15 downto 0) := (others => '0');
  signal pmul19_P2 :  std_logic_vector(15 downto 0) := (others => '0');
  signal pmul19_result :   std_logic_vector(15 downto 0);
  signal pmul19_tag_in: std_logic_vector(1 downto 0);
  signal pmul19_tag_out: std_logic_vector(1 downto 0);
  signal pmul19_start_req : std_logic := '0';
  signal pmul19_start_ack : std_logic := '0';
  signal pmul19_fin_req   : std_logic := '0';
  signal pmul19_fin_ack   : std_logic := '0';
  -- 
begin --
  -- clock/reset generation 
  clk <= not clk after 5 ns;
  -- assert reset for four clocks.
  process
  begin --
    Vhpi_Initialize;
    wait until clk = '1';
    wait until clk = '1';
    wait until clk = '1';
    wait until clk = '1';
    reset <= '0';
    while true loop --
      wait until clk = '0';
      Vhpi_Listen;
      Vhpi_Send;
      --
    end loop;
    wait;
    --
  end process;
  -- connect all the top-level modules to Vhpi
  process
  variable val_string, obj_ref: VhpiString;
  begin --
    wait until reset = '0';
    -- let the DUT come out of reset.... give it 4 cycles.
    wait until clk = '1';
    wait until clk = '1';
    wait until clk = '1';
    wait until clk = '1';
    while true loop -- 
      wait until clk = '0';
      wait for 1 ns;
      obj_ref := Pack_String_To_VHPI_String("pmul19 req");
      Vhpi_Get_Port_Value(obj_ref,val_string,1);
      pmul19_start_req <= To_Std_Logic(val_string);
      obj_ref := Pack_String_To_Vhpi_String("pmul19 0");
      Vhpi_Get_Port_Value(obj_ref,val_string, 16);
      pmul19_P1 <= Unpack_String(val_string,16);
      obj_ref := Pack_String_To_Vhpi_String("pmul19 1");
      Vhpi_Get_Port_Value(obj_ref,val_string, 16);
      pmul19_P2 <= Unpack_String(val_string,16);
      wait for 0 ns;
      if pmul19_start_req = '1' then -- 
        while true loop --
          wait until clk = '1';
          if pmul19_start_ack = '1' then exit; end if;--
        end loop; 
        pmul19_start_req <= '0';
        pmul19_fin_req <= '1';
        while true loop -- 
          wait until clk = '1';
          if pmul19_fin_ack = '1' then exit; end if; --  
        end loop; 
        pmul19_fin_req <= '0';
        -- 
      end if; 
      obj_ref := Pack_String_To_Vhpi_String("pmul19 ack");
      val_string := To_String(pmul19_fin_ack);
      Vhpi_Set_Port_Value(obj_ref,val_string,1);
      obj_ref := Pack_String_To_Vhpi_String("pmul19 0");
      val_string := Pack_SLV_To_Vhpi_String(pmul19_result);
      Vhpi_Set_Port_Value(obj_ref,val_string,16);
      -- 
    end loop;
    --
  end process;
  ahir_system_instance: ahir_system -- 
    port map ( -- 
      pmul19_P1 => pmul19_P1,
      pmul19_P2 => pmul19_P2,
      pmul19_result => pmul19_result,
      pmul19_tag_in => pmul19_tag_in,
      pmul19_tag_out => pmul19_tag_out,
      pmul19_start_req => pmul19_start_req,
      pmul19_start_ack => pmul19_start_ack,
      pmul19_fin_req  => pmul19_fin_req, 
      pmul19_fin_ack  => pmul19_fin_ack ,
      clk => clk,
      reset => reset); -- 
  -- 
end VhpiLink;
